library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library unisim;
use unisim.vcomponents.all;

entity Music5000_lx9core is
    port (
        -- System oscillator
        clk50        : in    std_logic;
        -- BBC 1MHZ Bus
        clke         : in    std_logic;
        rnw          : in    std_logic;
        rst_n        : in    std_logic;
        pgfc_n       : in    std_logic;
        pgfd_n       : in    std_logic;
        bus_addr     : in    std_logic_vector (7 downto 0);
        bus_data     : inout std_logic_vector (7 downto 0);
        bus_data_dir : out   std_logic;
        bus_data_oel : out   std_logic;
        nmi          : out   std_logic;
        irq          : out   std_logic;
        -- SPI DAC
        dac_cs_n     : out   std_logic;
        dac_sck      : out   std_logic;
        dac_sdi      : out   std_logic;
        dac_ldac_n   : out   std_logic;
        -- RAM (unused)
        ram_addr     : out   std_logic_vector(18 downto 0);
        ram_data     : inout std_logic_vector(7 downto 0);
        ram_cel      : out   std_logic;
        ram_oel      : out   std_logic;
        ram_wel      : out   std_logic;
        -- Misc
        pmod0        : out   std_logic_vector(7 downto 0);
        pmod1        : out   std_logic_vector(7 downto 0);
        pmod2        : in    std_logic_vector(3 downto 0);
        sw1          : in    std_logic;
        sw2          : in    std_logic;
        led          : out   std_logic
    );
end Music5000_lx9core;

architecture Behavioral of Music5000_lx9core is

signal clk6 : std_logic;
signal irq_n : std_logic;
signal spdif : std_logic;
signal filter : std_logic := '1';
signal sw1_out : std_logic := '0';
signal sw1_counter : unsigned(15 downto 0) := (others => '0');

begin

    ------------------------------------------------
    -- 6MHZ Clock Generation
    -- (from the 50.000MHZ Oscillator)
    ------------------------------------------------

    inst_DCM : DCM
        generic map (
            CLKFX_MULTIPLY   => 3,
            CLKFX_DIVIDE     => 25,
            CLKIN_PERIOD     => 20.000,
            CLK_FEEDBACK     => "NONE"
            )
        port map (
            CLKIN            => clk50,
            CLKFB            => '0',
            RST              => '0',
            DSSEN            => '0',
            PSINCDEC         => '0',
            PSEN             => '0',
            PSCLK            => '0',
            CLKFX            => clk6
            );

    ------------------------------------------------
    -- Music 5000 Core with SPI DAC Interface
    ------------------------------------------------

    inst_Music5000SpiDac : entity work.Music5000SpiDac
        generic map (
            sumwidth     => 19,
            dacwidth     => 18
            )
        port map (
            -- This is the 6MHz audio clock
            clk6         => clk6        ,
            -- This is the cpu clock
            clke         => clke        ,
            rnw          => rnw         ,
            rst_n        => rst_n       ,
            pgfc_n       => pgfc_n      ,
            pgfd_n       => pgfd_n      ,
            bus_addr     => bus_addr    ,
            bus_data     => bus_data    ,
            bus_data_oel => bus_data_oel,
            dac_cs_n     => dac_cs_n    ,
            dac_sck      => dac_sck     ,
            dac_sdi      => dac_sdi     ,
            dac_ldac_n   => dac_ldac_n  ,
            enable5      => '1'         ,
            enable3      => '1'         ,
            filter       => filter      ,
            spdif        => spdif       ,
            irq_n        => irq_n       ,
            owl          => pmod2(3)
            );

    ------------------------------------------------
    -- Filter off/on via sw1
    ------------------------------------------------
    process(clk6)
    begin
        if rising_edge(clk6) then
            if sw1 = sw1_out then
                sw1_counter <= (others => '0');
            else
                sw1_counter <= sw1_counter + 1;
                if sw1_counter = x"ffff" then
                    sw1_out <= sw1;
                    if sw1_out = '1' then
                        filter <= not filter;
                    end if;
                end if;
            end if;
        end if;
    end process;

    ------------------------------------------------
    -- 1MHZ Bus FPGA Adapter Specific Stuff
    ------------------------------------------------

    irq          <= not irq_n;
    nmi          <= '0';

    bus_data_dir <= rnw;

    ram_addr     <= (others => '0');
    ram_data     <= (others => '0');
    ram_cel      <= '1';
    ram_oel      <= '1';
    ram_wel      <= '1';

    pmod0        <= (others => '0');
    pmod1        <= "0" & spdif & "000000";

    led          <= filter;

end Behavioral;
